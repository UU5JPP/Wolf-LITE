
module DEBUG (
	probe);	

	input	[11:0]	probe;
endmodule
