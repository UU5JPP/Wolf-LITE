
module DEBUG2 (
	probe);	

	input	[23:0]	probe;
endmodule
